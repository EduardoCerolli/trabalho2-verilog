`timescale 1ns/1ps
module expandeChave_TB (
    
);
    
endmodule